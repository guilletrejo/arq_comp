`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
//	Alumnos:
//					 Ortmann, Nestor Javier
// 				 Trejo, Bruno Guillermo
// Year: 		 2018
// Module Name: MEMORIA DE DATOS
//////////////////////////////////////////////////////////////////////////////////
module DATA_MEM(
    );


endmodule
