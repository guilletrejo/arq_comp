`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// putarraqui
//////////////////////////////////////////////////////////////////////////////////
module MAIN(
    );
//soy nestor
// de una, soy guille
endmodule
