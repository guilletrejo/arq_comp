`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// putarraqui
//////////////////////////////////////////////////////////////////////////////////
module MAIN(
    );


endmodule
