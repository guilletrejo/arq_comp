`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
//	Alumnos:
//			     Ortmann, Nestor Javier
// 				 Trejo, Bruno Guillermo
// Year: 		 2019asdasda
// Module Name: TOP DI TUTTI TOPasdasdasd
//////////////////////////////////////////////////////////////////////////////////
module TOP(
    );


endmodule
