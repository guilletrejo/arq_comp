`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
//	Alumnos:
//					 Ortmann, Nestor Javier
// 				 Trejo, Bruno Guillermo
// Year: 		 2018
// Module Name: INSTRUCTION DECODER
//////////////////////////////////////////////////////////////////////////////////
module INSTRUCTION_DECODER(
    );


endmodule
