`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
//	Alumnos:
//					 Ortmann, Nestor Javier
// 				 Trejo, Bruno Guillermo
// Year: 		 2018
// Module Name: CONTROL
//////////////////////////////////////////////////////////////////////////////////
module CONTROL(
    );


endmodule
