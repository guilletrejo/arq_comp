`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
<<<<<<< HEAD
// Company: 
// Engineer: 
// 
// Create Date:    09:28:44 02/07/2019 
// Design Name: 
// Module Name:    REGISTERS 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module REGISTERS(
    );


endmodule
=======
//	Alumnos:
//				 Ortmann, Nestor Javier
// 				 Trejo, Bruno Guillermo
// Year: 		 2019
// Module Name:  REGISTROS
//////////////////////////////////////////////////////////////////////////////////

module REGISTERS#(
	parameter len_data = 32,
	parameter depth = 32,
	parameter num_bits = 5 //$clog2(depth)
	)
    (
	input clk,
	input reset,
	input RegWrite,
	input [num_bits-1:0] read_register_1,
	input [num_bits-1:0] read_register_2,
	input [num_bits-1:0] write_register,
	input [len_data-1:0] write_data,

	output [len_data-1:0] wire_read_data_1, // ver despues para que lo usa
	output reg [len_data-1:0] read_data_1,
	output reg [len_data-1:0] read_data_2
    );

	reg [len_data-1:0] registers_mips [depth-1:0]; // Banco de registros (tam. es len_data y cantidad es depth) 

	assign wire_read_data_1 = registers_mips[read_register_1]; // Algo desconozido aun

	generate
		integer i;		
		initial
        for (i = 0; i < depth; i = i + 1)
          registers_mips[i] = {len_data{1'b0+(i)}}; // reg0 = 0. reg1 = 1. reg2 = 2... etc.
	endgenerate

	always @(posedge clk)
	begin
		if (reset)
		begin
			read_data_1 <= 0;
			read_data_2 <= 0;
		end

		else begin
			read_data_1 <= registers_mips[read_register_1];
			read_data_2 <= registers_mips[read_register_2];
		end
	end

	always @(negedge clk)
	begin
		if (RegWrite) 
		begin
			registers_mips[write_register] <= write_data;				
		end
	end

endmodule
>>>>>>> 903dbfca61f1e992de6c9575a43a561051a84471
