`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
//	Alumnos:
//				 Ortmann, Nestor Javier
// 				 Trejo, Bruno Guillermo
// Year: 		 2019
// Module Name:  TOP MIPS
//////////////////////////////////////////////////////////////////////////////////

module TOP_MIPS#(
	parameter len_data = 32,
	parameter len_addr = 7,
	parameter len_test = 8,
	parameter num_bits = 5, //$clog2(len_data),
	parameter len_exec_bus = 11,
	parameter len_mem_bus = 9,
	parameter len_wb_bus = 2
	)(
	input clk,
	input reset,

	// para debug

	input debug_flag,
	input debug_ram_flag,
	input [len_data-1:0] debug_ram_addr,
	input [len_addr-1:0] in_addr_mem_inst,
	input [len_data-1:0] in_ins_to_mem,
	input wea_ram_inst,


	//PARA MANDAR A DEBUG.U
	output [len_data-1:0] out_reg0_recolector,
	output [len_data-1:0] out_reg1_recolector,
	output [len_data-1:0] out_reg2_recolector,
	output [len_data-1:0] out_reg3_recolector,
	output [len_data-1:0] out_reg4_recolector,
	output [len_data-1:0] out_reg5_recolector,
	output [len_data-1:0] out_reg6_recolector,
	output [len_data-1:0] out_reg7_recolector,
	output [len_data-1:0] out_pc,
	output [len_data-1:0] data0,
	output [len_data-1:0] data1,
	output [len_data-1:0] data2,
	output [len_data-1:0] data3,
	output [2*len_data-1:0] Latch_IF_ID,
	output [4*len_data-1:0] Latch_ID_EX,
	output [4*len_data-1:0] Latch_EX_MEM,
	output [3*len_data-1:0] Latch_MEM_WB,
	//----------------------------------------

	output [len_test-1:0] out_inst_test,
	output halt_flag
	);

    wire [len_data-1:0] connect_in_pc_branch_1_2,
				   connect_in_pc_branch_2_3,
				   connect_in_pc_jump,
				   connect_in_pc_jump_register,
				   connect_instruccion,
				   connect_reg1,
				   connect_reg2,
				   connect_sign_extend,
				   connect_alu_out,
				   connect_write_data_5_2,
				   connect_read_data,
				   connect_out_addr_mem,
				   connect_write_data_3_4,
				   connect_in_pc_branch_3_4,
				   connect_in_pc_branch_4_1,
				   connect_reg0_recolector,
				   connect_reg1_recolector,
				   connect_reg2_recolector,
				   connect_reg3_recolector,
				   connect_reg4_recolector,
				   connect_reg5_recolector,
				   connect_reg6_recolector,
				   connect_reg7_recolector,
				   connect_out_pc,
				   out_data_debug;
	wire [len_test-1:0] conn_inst_test; // va a los led

	wire [num_bits-1:0] connect_rt,
						connect_rd,
						connect_rs,
						connect_shamt,
						connect_write_reg_3_4,
						connect_write_reg_4_2;

    wire [len_exec_bus-1:0] connect_execute_bus;
	
	wire [len_mem_bus-1:0] connect_memory_bus_2_3,
			   connect_memory_bus_3_4;
	
	wire [len_wb_bus-1:0] connect_writeBack_bus_2_3,
			   connect_out_writeBack_bus,
			   connect_writeBack_bus_3_4;
    
    wire connect_flag_jump,
         connect_flag_jump_register,
	     connect_zero_flag,
	     connect_branch_flag,
	     connect_stall_flag,
	     connect_halt_flag_1_2,
	     connect_halt_flag_2_3,
	     connect_halt_flag_3_4,
	     connect_halt_flag_4_5; 

	assign connect_write_data_5_2 = (connect_out_writeBack_bus[0]) ? connect_read_data : connect_out_addr_mem;

	/* Para mandar a Debug Unit */
	assign out_reg0_recolector = connect_reg0_recolector;
	assign out_reg1_recolector = connect_reg1_recolector;
	assign out_reg2_recolector = connect_reg2_recolector;
	assign out_reg3_recolector = connect_reg3_recolector;
	assign out_reg4_recolector = connect_reg4_recolector;
	assign out_reg5_recolector = connect_reg5_recolector;
	assign out_reg6_recolector = connect_reg6_recolector;
	assign out_reg7_recolector = connect_reg7_recolector;
	assign out_pc = connect_out_pc;
	assign data0 = out_data_debug;
	assign data1 = out_data_debug;
	assign data2 = out_data_debug;
	assign data3 = out_data_debug;
	
	assign Latch_IF_ID = {	// 2 registros TOTAL 64 BITS
		connect_instruccion, // 32 bits
		connect_in_pc_branch_1_2 // 32 bits
	};
	assign Latch_ID_EX = {	// 4 registros 		TOTAL 128 BITS
		{10{1'b 0}}, // 10 bits --> Se agrega para alinear
		connect_execute_bus, // 11 bits
		connect_memory_bus_2_3, // 9 bits
		connect_writeBack_bus_2_3, // 2 bits
		{12{1'b 0}}, // 12 bits --> Se agrega para alinear
		connect_rd, // 5 bits
		connect_rs, // 5 bits
		connect_rt, // 5 bits
		connect_shamt, // 5 bits
		connect_sign_extend, // 32 bits
		connect_in_pc_branch_2_3 // 32 bits
	};
	assign Latch_EX_MEM = {	// 4 registros		TOTAL 128 BITS
		{15{1'b 0}}, // 15 bits
		connect_memory_bus_3_4, // 9 bits
		connect_writeBack_bus_3_4, // 2 bits
		connect_write_reg_3_4, // 5 bits
		connect_zero_flag, // 1 bit
		connect_alu_out, // 32 bits
		connect_in_pc_branch_3_4, // 32 bits
		connect_reg1 // 32 bits
	};

	assign Latch_MEM_WB = {	// 4 registros 		TOTAL 128 BITS
		{24{1'b 0}}, // 24 bits
		connect_halt_flag_4_5, // 1 bitconnect_stall_flag
		connect_write_reg_4_2, // 5 bits
		connect_out_writeBack_bus, // 2 bits
		connect_out_addr_mem, // 32 bits
		connect_read_data // 32 bits
	};
	/* ------------------------ */
	
	assign out_inst_test = conn_inst_test;
	assign halt_flag = connect_halt_flag_4_5;

	IF_ID #(
		.len_data(len_data)
		)
		u_if_id(
			.clk(clk),
			.reset(reset),
			.in_pc_src({connect_flag_jump, connect_flag_jump_register, connect_branch_flag}),
			.in_pc_jump(connect_in_pc_jump),
			.in_branch_address(connect_in_pc_branch_4_1),
			.in_pc_register(connect_in_pc_jump_register),
			.stall_flag(connect_stall_flag),

			.in_addr_debug(in_addr_mem_inst),
			.debug_flag(debug_flag),
			.in_ins_to_mem(in_ins_to_mem),
			.wea_ram_inst(wea_ram_inst),

			.out_pc_branch(connect_in_pc_branch_1_2),
			.out_instruction(connect_instruccion),
			.out_pc(connect_out_pc), 
			.out_inst_test(conn_inst_test),
			.out_halt_flag_if(connect_halt_flag_1_2) 
		);

	ID_EX #(
		.len_data(len_data)
		)
		u_id_ex(
			.clk(clk),
			.reset(reset),
			.in_pc_branch(connect_in_pc_branch_1_2),
			.in_instruccion(connect_instruccion),

			.RegWrite(connect_out_writeBack_bus[1]),
			.write_data(connect_write_data_5_2),
			.write_register(connect_write_reg_4_2),
			.flush(connect_branch_flag),
			
			.out_pc_branch(connect_in_pc_branch_2_3),
			.out_pc_jump(connect_in_pc_jump),
			.out_pc_jump_register(connect_in_pc_jump_register),
			.out_reg1(connect_reg1),
			.out_reg2(connect_reg2),
			.out_sign_extend(connect_sign_extend),
			.out_rt(connect_rt),
			.out_rd(connect_rd),
			.out_rs(connect_rs),
			.out_shamt(connect_shamt),

			.out_reg0_recolector(connect_reg0_recolector),
			.out_reg1_recolector(connect_reg1_recolector),
			.out_reg2_recolector(connect_reg2_recolector),
			.out_reg3_recolector(connect_reg3_recolector),
			.out_reg4_recolector(connect_reg4_recolector),
			.out_reg5_recolector(connect_reg5_recolector),
			.out_reg6_recolector(connect_reg6_recolector),
			.out_reg7_recolector(connect_reg7_recolector),

			.execute_bus(connect_execute_bus),
			.flag_jump(connect_flag_jump),
			.flag_jump_register(connect_flag_jump_register),
			.memory_bus(connect_memory_bus_2_3),
			.writeBack_bus(connect_writeBack_bus_2_3),

			.stall_flag(connect_stall_flag),

			.halt_flag_d(connect_halt_flag_1_2),
			.out_halt_flag_d(connect_halt_flag_2_3)
		);

	EX_MEM #(
		.len_data(len_data)
		)
		u_ex_mem(
			.clk(clk),
			.reset(reset),
		
			.in_pc_branch(connect_in_pc_branch_2_3),
			.in_reg1(connect_reg1),
			.in_reg2(connect_reg2),
			.in_sign_extend(connect_sign_extend),
			.in_rt(connect_rt),
			.in_rd(connect_rd),
			.in_shamt(connect_shamt),
		
			.execute_bus(connect_execute_bus),
			.memory_bus(connect_memory_bus_2_3),
			.writeBack_bus(connect_writeBack_bus_2_3), 

			.ex_mem_reg_write(connect_writeBack_bus_3_4[1]),
			.mem_wb_reg_write(connect_out_writeBack_bus[1]),
			.ex_mem_rd(connect_write_reg_3_4),
			.mem_wb_rd(connect_write_reg_4_2),
			.in_rs(connect_rs),

			.in_mem_forw(connect_alu_out),
			.in_wb_forw(connect_write_data_5_2),
			.flush(connect_branch_flag),
		
			.out_pc_branch(connect_in_pc_branch_3_4),
			.out_alu(connect_alu_out),
			.zero_flag(connect_zero_flag),
			.out_reg2(connect_write_data_3_4),
			.out_write_reg(connect_write_reg_3_4),
		
			// señales de control
			.memory_bus_out(connect_memory_bus_3_4),
			.writeBack_bus_out(connect_writeBack_bus_3_4),

			.halt_flag_e(connect_halt_flag_2_3),
			.out_halt_flag_e(connect_halt_flag_3_4)
			);

	MEM_WB #(
		.len_data(len_data)
		)
		u_mem_wb(
			.clk(clk),
			.reset(reset),
			.in_addr_mem(debug_ram_flag? debug_ram_addr : connect_alu_out),
			.write_data(connect_write_data_3_4),
			
			.memory_bus(connect_memory_bus_3_4),
		    .in_writeBack_bus(connect_writeBack_bus_3_4),
			.in_write_reg(connect_write_reg_3_4),			
			.zero_flag(connect_zero_flag),
			.in_pc_branch(connect_in_pc_branch_3_4),
			.halt_flag_m(connect_halt_flag_3_4),

			//outputs		
			.read_data(connect_read_data),
			.pc_src(connect_branch_flag),
			.out_pc_branch(connect_in_pc_branch_4_1),
		    .out_writeBack_bus(connect_out_writeBack_bus),
			.out_addr_mem(connect_out_addr_mem),
			.out_write_reg(connect_write_reg_4_2),

			//para mostrar en debug unit
			.out_data_debug(out_data_debug),
			//

			.out_halt_flag_m(connect_halt_flag_4_5)
			);

endmodule
